module segment_7 (in, HEX);
   input [3:0] in;
	output [0:6] HEX;
	assign HEX=(in==4'b0000) ? 7'b0000001:
	           (in==4'b0001) ? 7'b1001111:
	           (in==4'b0010) ? 7'b0010010:
				  (in==4'b0011) ? 7'b0000110:
				  (in==4'b0100) ? 7'b1001100:
				  (in==4'b0101) ? 7'b0100100:
				  (in==4'b0110) ? 7'b0100000:
				  (in==4'b0111) ? 7'b0001101:
				  (in==4'b1000) ? 7'b0000000:
				  (in==4'b1001) ? 7'b0000100:
                              7'b1111111;
endmodule